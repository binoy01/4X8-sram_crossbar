module ad3(input [8:0] a3, input [10:0] b3, output reg [11:0] c3
    );



always@(*)

c3= a3+b3;
    
endmodule
