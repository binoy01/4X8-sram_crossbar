module mult(input [3:0] a, input [3:0] b, output reg [8:0] c
    );

always@(*)

c= a*b;


endmodule
