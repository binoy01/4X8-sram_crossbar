module ad2(input [8:0] a2, input [9:0] b2, output reg [10:0] c2
    );



always@(*)

c2= a2+b2;
