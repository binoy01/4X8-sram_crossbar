module ad(input [8:0] a1, input [8:0] b1, output reg [9:0] c1
    );



always@(*)

c1= a1+b1;
    
   
endmodule
